** Generated for: hspiceD
** Generated on: Sep 12 18:42:00 2023
** Design library name: test
** Design cell name: inverter
** Design view name: schematic




** Library name: test
** Cell name: inverter
** View name: schematic
m0 y a vss vss nmos_rvt w=81e-9 l=20e-9 nfin=3
m1 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
.END
